`timescale 1ns / 1ps

module ComparatorTb();
    reg  [2:0] q;
    reg  [1:0] s;
    wire [2:0] result;
    
    Comparator uut(
        .q(q),
        .s(s),
        .result(result)
    );
    
    initial begin
        q = 0; s = 0;
        #100;
        q = 0; s = 1;
        #100;
        q = 0; s = 2;
        #100;
        q = 0; s = 3;
        #100;
        q = 1; s = 0;
        #100;
        q = 1; s = 1;
        #100;
        q = 1; s = 2;
        #100;
        q = 1; s = 3;
        #100;
        q = 2; s = 0;
        #100;
        q = 2; s = 1;
        #100;
        q = 2; s = 2;
        #100;
        q = 2; s = 3;
        #100;
        
        q = 3; s = 0;
        #100;
        q = 3; s = 1;
        #100;
        q = 3; s = 2;
        #100;
        q = 3; s = 3;
        #100;
        q = 4; s = 0;
        #100;
        q = 4; s = 1;
        #100;
        q = 4; s = 2;
        #100;
        q = 4; s = 3;
        #100;
        q = 5; s = 0;
        #100;
        q = 5; s = 1;
        #100;
        q = 5; s = 2;
        #100;
        q = 5; s = 3;
        #100;
        
        q = 6; s = 0;
        #100;
        q = 6; s = 1;
        #100;
        q = 6; s = 2;
        #100;
        q = 6; s = 3;
        #100;
        q = 7; s = 0;
        #100;
        q = 7; s = 1;
        #100;
        q = 7; s = 2;
        #100;
        q = 7; s = 3;
        #100;
        
    end
endmodule